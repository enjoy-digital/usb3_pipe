parameter	[7:0]	DESCR_USB2_DEVICE	= 'd0;
parameter	[6:0]	DESCR_USB3_DEVICE	= 'd0;
parameter	[7:0]	DESCR_USB2_DEVICE_QUAL	= 'd18;
parameter	[7:0]	DESCR_USB2_CONFIG	= 'd28;
parameter	[6:0]	DESCR_USB3_CONFIG	= 'd5;
parameter	[7:0]	DESCR_USB2_CONFIG_LEN	= 'd41;
parameter	[6:0]	DESCR_USB3_CONFIG_LEN	= 'd53;
parameter	[6:0]	DESCR_USB3_BOS    	= 'd19;
parameter	[6:0]	DESCR_USB3_BOS_LEN	= 'd22;
parameter	[7:0]	DESCR_USB2_STRING0	= 'd69;
parameter	[6:0]	DESCR_USB3_STRING0	= 'd25;
parameter	[7:0]	DESCR_USB2_STRING1	= 'd73;
parameter	[6:0]	DESCR_USB3_STRING1	= 'd26;
parameter	[7:0]	DESCR_USB2_STRING2	= 'd113;
parameter	[6:0]	DESCR_USB3_STRING2	= 'd36;
parameter	[7:0]	DESCR_USB2_STRING3	= 'd145;
parameter	[6:0]	DESCR_USB3_STRING3	= 'd44;
parameter	[7:0]	DESCR_USB2_CONFUNSET	= 'd171;
parameter	[6:0]	DESCR_USB3_CONFUNSET	= 'd51;
parameter	[7:0]	DESCR_USB2_CONFSET	= 'd172;
parameter	[6:0]	DESCR_USB3_CONFSET	= 'd52;
parameter	[7:0]	DESCR_USB2_EOF     	= 'd173;
parameter	[6:0]	DESCR_USB3_EOF     	= 'd53;
