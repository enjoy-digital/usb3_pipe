parameter	[7:0]	DESCR_USB2_DEVICE	= 'd0;
parameter	[6:0]	DESCR_USB3_DEVICE	= 'd0;
parameter	[7:0]	DESCR_USB2_DEVICE_QUAL	= 'd0;
parameter	[7:0]	DESCR_USB2_CONFIG	= 'd0;
parameter	[6:0]	DESCR_USB3_CONFIG	= 'd0;
parameter	[7:0]	DESCR_USB2_CONFIG_LEN	= 'd41;
parameter	[6:0]	DESCR_USB3_CONFIG_LEN	= 'd53;
parameter	[6:0]	DESCR_USB3_BOS    	= 'd0;
parameter	[6:0]	DESCR_USB3_BOS_LEN	= 'd22;
parameter	[7:0]	DESCR_USB2_STRING0	= 'd0;
parameter	[6:0]	DESCR_USB3_STRING0	= 'd0;
parameter	[7:0]	DESCR_USB2_STRING1	= 'd0;
parameter	[6:0]	DESCR_USB3_STRING1	= 'd0;
parameter	[7:0]	DESCR_USB2_STRING2	= 'd0;
parameter	[6:0]	DESCR_USB3_STRING2	= 'd0;
parameter	[7:0]	DESCR_USB2_STRING3	= 'd0;
parameter	[6:0]	DESCR_USB3_STRING3	= 'd0;
parameter	[7:0]	DESCR_USB2_CONFUNSET	= 'd0;
parameter	[6:0]	DESCR_USB3_CONFUNSET	= 'd0;
parameter	[7:0]	DESCR_USB2_CONFSET	= 'd0;
parameter	[6:0]	DESCR_USB3_CONFSET	= 'd0;
parameter	[7:0]	DESCR_USB2_EOF     	= 'd0;
parameter	[6:0]	DESCR_USB3_EOF     	= 'd0;
